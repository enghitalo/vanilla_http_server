module http1_1
