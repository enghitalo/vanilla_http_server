module http2

// HPACK header compression/decompression stubs (RFC 7541)
// TODO: Implement full HPACK encoder/decoder

pub struct HpackDecoder {}

pub struct HpackEncoder {}
